module top_module ( input a, input b, output out );
    mod_a left_side (a,b,out );
endmodule
